module vga_pic(
	input wire vga_clk,
	input wire sys_rst_n,
	input wire [9:0] pix_x,
	input wire [9:0] pix_y,
	output reg [15:0] pix_data
);

parameter   CHAR_B_H = 10'd140,
            CHAR_B_V = 10'd216,
				CHAR_W = 10'd256,
            CHAR_H = 10'd128,
            BLACK = 16'h0000,
            WHITE = 16'hFFFF,
            GOLDEN = 16'hFEC0;

wire [9:0] char_x;
wire [9:0] char_y;

reg [255:0] char [127:0];

assign  char_x  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_x - CHAR_B_H) : 10'h3FF;
assign  char_y  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_y - CHAR_B_V) : 10'h3FF;

always@(posedge vga_clk)
    begin
        char[0]     <=  256'h00000000000000000000000000000000;
        char[1]     <=  256'h00000000000000000000000000000000;
        char[2]     <=  256'h00000000000000000000000000000000;
        char[3]     <=  256'h00000000000000000000000000000000;
        char[4]     <=  256'h00000000000000000000000000000000;
        char[5]     <=  256'h00000000000000000000000000000000;
        char[6]     <=  256'h00000000000000000000000000000000;
        char[7]     <=  256'h00000000000000000000000000000000;
        char[8]     <=  256'h00000000000000000000000000000000;
        char[9]     <=  256'h00000000000000000000000000000000;
        char[10]    <=  256'h00000000000000000000000000000000;
        char[11]    <=  256'hFF8003FF7FF807FE001FE0000FFFFFF0;
        char[12]    <=  256'hFF8003FF7FF807FE007FF8800FFFFFF0;
        char[13]    <=  256'h1F8003F80FC000F000F03F800F03C0F8;
        char[14]    <=  256'h1F8003F80780006001C00F801E03C038;
        char[15]    <=  256'h1F8007F80780006003C007801C03C038;
        char[16]    <=  256'h1FC007F807800060078003C01803C018;
        char[17]    <=  256'h1FC007F807800060078001C01803C018;
        char[18]    <=  256'h1FC007F807800060070001C01003C00C;
        char[19]    <=  256'h1FC00FF8078000600F0000C03003C00C;
        char[20]    <=  256'h1FE00FF8078000600F0000C03003C004;
        char[21]    <=  256'h1FE00FF8078000600F0000000003C000;
        char[22]    <=  256'h1FE00FF8078000600F0000000003C000;
        char[23]    <=  256'h1FE00FF8078000600F0000000003C000;
        char[24]    <=  256'h1FE01FF8078000600F8000000003C000;
        char[25]    <=  256'h1FF01FF80780006007C000000003C000;
        char[26]    <=  256'h1FF01DF80780006007E000000003C000;
        char[27]    <=  256'h1DF01DF80780006007F000000003C000;
        char[28]    <=  256'h1DF03DF80780006003FC00000003C000;
        char[29]    <=  256'h1DF83DF80780006001FF00000003C000;
        char[30]    <=  256'h1DF839F807800060007FC0000003C000;
        char[31]    <=  256'h1CF839F807800060003FF0000003C000;
        char[32]    <=  256'h1CF879F807800060000FFC000003C000;
        char[33]    <=  256'h1CF879F8078000600003FE000003C000;
        char[34]    <=  256'h1CFC71F8078000600000FF000003C000;
        char[35]    <=  256'h1C7C71F80780006000003F800003C000;
        char[36]    <=  256'h1C7CF1F80780006000000FC00003C000;
        char[37]    <=  256'h1C7CF1F807800060000007E00003C000;
        char[38]    <=  256'h1C7EE1F807800060000003E00003C000;
        char[39]    <=  256'h1C7EE1F807800060000001E00003C000;
        char[40]    <=  256'h1C3EE1F807800060000001F00003C000;
        char[41]    <=  256'h1C3FE1F807800060000000F00003C000;
        char[42]    <=  256'h1C3FE1F807800060080000F00003C000;
        char[43]    <=  256'h1C3FC1F807800060180000F00003C000;
        char[44]    <=  256'h1C1FC1F807800060180000F00003C000;
        char[45]    <=  256'h1C1FC1F8078000601C0000F00003C000;
        char[46]    <=  256'h1C1FC1F8078000600C0000F00003C000;
        char[47]    <=  256'h1C1F81F8078000E00E0000E00003C000;
        char[48]    <=  256'h1C1F81F8038000C00E0001E00003C000;
        char[49]    <=  256'h1C0F81F803C001C00F0001C00003C000;
        char[50]    <=  256'h1C0F81F801C003800F8003C00003C000;
        char[51]    <=  256'h1C0F01F801E007000FC007800003C000;
        char[52]    <=  256'hFF8F0FFF00F81E0007F81F000007E000;
        char[53]    <=  256'hFF870FFF003FFC00061FFC00007FFE00;
        char[54]    <=  256'h00000000000FE0000407F000007FFE00;
        char[55]    <=  256'h00000000000000000000000000000000;
        char[56]    <=  256'h00000000000000000000000000000000;
        char[57]    <=  256'h00000000000000000000000000000000;
        char[58]    <=  256'h00000000000000000000000000000000;
        char[59]    <=  256'h00000000000000000000000000000000;
        char[60]    <=  256'h00000000000000000000000000000000;
        char[61]    <=  256'h00000000000000000000000000000000;
        char[62]    <=  256'h00000000000000000000000000000000;
        char[63]    <=  256'h00000000000000000000000000000000;	  
    end

always@(posedge vga_clk or negedge sys_rst_n)
    if(sys_rst_n == 1'b0)
        pix_data    <= BLACK;
    else    if((((pix_x >= (CHAR_B_H - 1'b1))
                && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
                && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                && (char[char_y][10'd255 - char_x] == 1'b1))
        pix_data    <=  GOLDEN;
    else
        pix_data    <=  BLACK;

endmodule
